module CommTB()




endmodule

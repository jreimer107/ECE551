module CommTB();




endmodule
